.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt OAI21 Y A B1 B2
 XN1 A 0 intN RV523_NMOS
 XN2 B1 intN Y RV523_NMOS
 XN3 B2 intN Y RV523_NMOS
 XP1 A VDD Y RV523_PMOS
 XP2 B1 VDD intB RV523_PMOS
 XP3 B2 intB Y RV523_PMOS
.ends
