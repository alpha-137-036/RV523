module BUF(
    output Y,
    input A
);
    assign Y = A;
endmodule