.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt NOR3 Y A B C
 XN1 A 0 Y RV523_NMOS
 XN2 B 0 Y RV523_NMOS
 XN3 C 0 Y RV523_NMOS
 XP1 A int1 Y RV523_PMOS
 XP2 B int2 int1 RV523_PMOS
 XP3 C VDD int2 RV523_PMOS
.ends
