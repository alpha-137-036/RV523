module DECAP();
endmodule