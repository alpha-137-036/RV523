.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt NOR Y A B
 XN1 A 0 Y RV523_NMOS
 XN2 B 0 Y RV523_NMOS
 XP1 A VDD C RV523_PMOS
 XP2 B C Y RV523_PMOS
.ends
