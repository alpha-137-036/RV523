.subckt NOR3 Y A1 A2 A3 VDD VSS
 XN1 A1 VSS Y RV523_NMOS
 XN2 A2 VSS Y RV523_NMOS
 XN3 A3 VSS Y RV523_NMOS
 XP1 A1 int1 Y RV523_PMOS
 XP2 A2 int2 int1 RV523_PMOS
 XP3 A3 VDD int2 RV523_PMOS
.ends
