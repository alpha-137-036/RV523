.subckt NAND3 A B C Y
X0 int1 A 0 N7002
X1 int2 B int1 N7002
X2 Y C int2 N7002
X3 Y A VDD BSS84
X4 Y B VDD BSS84
X5 Y C VDD BSS84
.ends


