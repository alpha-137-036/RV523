.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt AOI211 Y A B C1 C2
 XN1 A 0 Y RV523_NMOS
 XN2 B 0 Y RV523_NMOS
 XN3 C1 0 intC RV523_NMOS
 XN4 C2 intC Y RV523_NMOS
 XP1 A VDD intPA RV523_PMOS
 XP2 B intPA intPB RV523_PMOS
 XP3 C1 intPB Y RV523_PMOS
 XP4 C2 intPB Y RV523_PMOS
.ends
