* Main ngspice simulation file

.include "../RV523_global.sp"
.include "OAI211.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A B C1 C2 VDD 0 OAI211

.TRAN 0.1ns 48200ns

* Simulation control
.control 
    run
    write OAI211.raw
    quit
.endc
.END