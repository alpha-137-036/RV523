module AND2(
    output Y,
    input A1,
    input A2
);
    assign Y = A1 & A2;
endmodule