.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt OAI22 Y A1 A2 B1 B2
 XN1 A1 0 intN RV523_NMOS
 XN2 A2 0 intN RV523_NMOS
 XN3 B1 intN Y RV523_NMOS
 XN4 B2 intN Y RV523_NMOS
 XP1 A1 VDD intA RV523_PMOS
 XP2 A2 intA Y RV523_PMOS
 XP3 B1 VDD intB RV523_PMOS
 XP4 B2 intB Y RV523_PMOS
.ends
