* Main ngspice simulation file

.include "NAND3.ckt"
.include "pwl_Inputs.sp"
.include "../2n7002.sub"
.include "../bss84.sub"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate NAND gate
XU1 A B C Y NAND3

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write NAND3.raw
    quit
.endc
.END