.subckt SR_LATCH Q nQ nS nR VDD VSS
 XN1 nS VSS intN1 RV523_NMOS
 XN2 nQ intN1 Q RV523_NMOS
 XN3 nR VSS intN2 RV523_NMOS
 XN4 Q intN2 nQ RV523_NMOS
 XP1 nS VDD Q RV523_PMOS
 XP2 nQ VDD Q RV523_PMOS
 XP3 nR VDD nQ RV523_PMOS
 XP4 Q VDD nQ RV523_PMOS
.ends
