.subckt NOR2 Y A1 A2 VDD VSS
 XN1 A1 VSS Y RV523_NMOS
 XN2 A2 VSS Y RV523_NMOS
 XP1 A1 VDD C RV523_PMOS
 XP2 A2 C Y RV523_PMOS
.ends
