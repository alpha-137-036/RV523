module NAND4(
    output Y,
    input A1,
    input A2,
    input A3,
    input A4
);
    assign Y = ~(A1 & A2 & A3 & A4);
endmodule