module NOT(
    output Y,
    input A
);
    assign Y = !A;
endmodule