* Main ngspice simulation file

.include "NOR3.ckt"
.include "pwl_Inputs.sp"
.include "../2n7002.sub"
.include "../bss84.sub"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate cell
XU1 A B C Y NOR3

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write NOR3.raw
    quit
.endc
.END