.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt NOR4 Y A1 A2 A3 A4
 XN1 A1 0 Y RV523_NMOS
 XN2 A2 0 Y RV523_NMOS
 XN3 A3 0 Y RV523_NMOS
 XN4 A4 0 Y RV523_NMOS
 XP1 A1 int1 Y RV523_PMOS
 XP2 A2 int2 int1 RV523_PMOS
 XP3 A3 int3 int2 RV523_PMOS
 XP4 A4 VDD int3 RV523_PMOS
.ends
