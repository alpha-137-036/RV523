.subckt BUF Y A VDD VSS
 Xnot1.N1 A VSS nA RV523_NMOS
 Xnot1.P1 A VDD nA RV523_PMOS
 Xnot2.N1 nA VSS Y RV523_NMOS
 Xnot2.P1 nA VDD Y RV523_PMOS
.ends
