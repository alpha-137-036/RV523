* Main ngspice simulation file

.include "NOR3.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate cell
XU1 Y A1 A2 A3 NOR3

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write NOR3.raw
    quit
.endc
.END