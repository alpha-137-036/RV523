* Main ngspice simulation file

.include "../RV523_global.sp"
.include "OAI21.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A B1 B2 VDD 0 OAI21

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write OAI21.raw
    quit
.endc
.END