* Main ngspice simulation file

.include "../RV523_global.sp"
.include "NAND3.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate NAND gate
XU1 Y A1 A2 A3 VDD 0 NAND3

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write NAND3.raw
    quit
.endc
.END