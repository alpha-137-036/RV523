* file alu.cir

.include 2n7002.sub
.include bss84.sub

* the power supply 3.3 V
Vcc cc0 0 3.3
Rcc cc cc0 10

Cdec 0 cc 10u

.global cc

.SUBCKT NOT A Y

XNnA Y A 0 N7002
XPnA Y A cc BSS84
.ENDS XOR

.SUBCKT NAND A B Y 

XPA Y A cc BSS84
XPB Y B cc BSS84

XNA Y A x1 N7002
XNB x1 B 0 N7002
.ENDS NAND

.SUBCKT AND A B Y
Xnand A B nY NAND
Xinv nY Y NOT
.ENDS AND

.SUBCKT NOR A B Y
XPA Y A p1 BSS84
XPB p1 B cc BSS84

XNA Y A 0 N7002
XNB Y B 0 N7002

.ENDS NOR

.SUBCKT OR A B Y
Xnor A B nY NOR
Xinv nY Y NOT
.ENDS OR

.SUBCKT AOI22 A1 A2 B1 B2 Y

XN1 xn1 A1 0 N7002
XN2 Y A2 xn1 N7002
XN3 xn2 B1 0 N7002
XN4 Y B2 xn2 N7002

XP1 Y B1 xp BSS84
XP2 Y B2 xp BSS84
XP3 xp A1 cc BSS84
XP4 xp A2 cc BSS84

.ENDS AOI22

.SUBCKT XOR A B Y

XnA A nA NOT
XnB B nB NOT

Xx A B nA nB Y AOI22
.ENDS XOR

.SUBCKT SLICE SUB nSUB A B nG P 

XnA A nA NOT

Xx A SUB nA nSUB AxSUB AOI22

XnG AxSUB B nG NAND
XP AxSUB B P OR

.ENDS SLICE 

Xslice0 SUB nSUB A0 B0 nG0 P0 SLICE
Xslice1 SUB nSUB A1 B1 nG1 P1 SLICE
Xslice2 SUB nSUB A2 B2 nG2 P2 SLICE
Xslice3 SUB nSUB A3 B3 nG3 P3 SLICE
Xslice4 SUB nSUB A4 B4 nG4 P4 SLICE
Xslice5 SUB nSUB A5 B5 nG5 P5 SLICE
Xslice6 SUB nSUB A6 B6 nG6 P6 SLICE
Xslice7 SUB nSUB A7 B7 nG7 P7 SLICE

.SUBCKT CLAH nG1 P1 nG2 P2 nG 
XG1 nG1 nG2 x1 NAND
XG2 x1 P2 nG NAND
.ENDS CLA

.SUBCKT CLA nG1 P1 nG2 P2 nG P 
XG1 nG1 nG2 x1 NAND
XG2 x1 P2 nG NAND
XP1 P1 P2 x2 NAND
XP2 x2 nG P NAND
.ENDS CLA

XCLA10 nG0 P0 nG1 P1 nG10 P10 CLA
XCLA32 nG2 P2 nG3 P3 nG32 P32 CLA
XCLA54 nG4 P4 nG5 P5 nG54 P54 CLA
XCLA76 nG6 P6 nG7 P7 nG76 P76 CLA

XCLA30 nG10 P10 nG32 P32 nG30 P30 CLA
XCLA74 nG54 P54 nG76 P76 nG74 P74 CLA

XCLA70 nG30 P30 nG74 P74 nG70 CLAH

XCLA20 nG10 P10 nG2 P2 nG20 P20 CLA

XCLA40 nG30 P30 nG4 P4 nG40 P40 CLA
XCLA50 nG30 P30 nG54 P54 nG50 P50 CLA

XCLA64 nG54 P54 nG6 P6 nG64 P64 CLA
XCLA60 nG30 P30 nG64 P64 nG60 P60 CLA


* the input signal for dc and tran simulation
aIn 
+ [DSUB DnSUB DA0 DA1 DA2 DA3 DA4 DA5 DA6 DA7 DB0 DB1 DB2 DB3 DB4 DB5 DB6 DB7] input_vector
 .model input_vector d_source(input_file = "alu_test_vectors.txt")

aInBridge 
+[DSUB DnSUB DA0 DA1 DA2 DA3 DA4 DA5 DA6 DA7 DB0 DB1 DB2 DB3 DB4 DB5 DB6 DB7]
+[SUB nSUB A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7] dac1
.model dac1 dac_bridge(out_low=0 out_high=3.3 out_undef=2.2 t_rise=10e-9 t_fall=10e-9  input_load = 5.0e-12)

aOutBridge 
+[nG70 nG60] 
+[DnG70 DnG60] adc1
.model adc1 adc_bridge(in_low=1 in_high=2)

* simulation commands
.tran 1n 20u

.control
    run
    write alu.raw cc I(Vcc) nG60 nG70
    eprvcd DSUB DnSUB DA0 DA1 DA2 DA3 DA4 DA5 DA6 DA7 DB0 DB1 DB2 DB3 DB4 DB5 DB6 DB7 DnG60 DnG70 > alu_out.vcd
.endc

.end