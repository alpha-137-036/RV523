.subckt AOI211 Y A B C1 C2 VDD VSS
 XN1 A VSS Y RV523_NMOS
 XN2 B VSS Y RV523_NMOS
 XN3 C1 VSS intC RV523_NMOS
 XN4 C2 intC Y RV523_NMOS
 XP1 A VDD intPA RV523_PMOS
 XP2 B intPA intPB RV523_PMOS
 XP3 C1 intPB Y RV523_PMOS
 XP4 C2 intPB Y RV523_PMOS
.ends
