module XNOR2(
    output Y,
    input A,
    input B
);
    assign Y = ~(A ^ B);
endmodule