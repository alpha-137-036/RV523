.subckt XOR2 Y A B VDD VSS
 Xaoi.N1 A VSS aoi.intA RV523_NMOS
 Xaoi.N2 B aoi.intA Y RV523_NMOS
 Xaoi.N3 aoi.B1 VSS aoi.intB RV523_NMOS
 Xaoi.N4 aoi.B2 aoi.intB Y RV523_NMOS
 Xaoi.P1 A aoi.intP Y RV523_PMOS
 Xaoi.P2 B aoi.intP Y RV523_PMOS
 Xaoi.P3 aoi.B1 VDD aoi.intP RV523_PMOS
 Xaoi.P4 aoi.B2 VDD aoi.intP RV523_PMOS
 XnotA.N1 A VSS aoi.B1 RV523_NMOS
 XnotA.P1 A VDD aoi.B1 RV523_PMOS
 XnotB.N1 B VSS aoi.B2 RV523_NMOS
 XnotB.P1 B VDD aoi.B2 RV523_PMOS
.ends
