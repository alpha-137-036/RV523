.subckt NOT Y A VDD VSS
 XN1 A VSS Y RV523_NMOS
 XP1 A VDD Y RV523_PMOS
.ends
