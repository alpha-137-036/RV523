.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt SR_LATCH Q nQ nS nR
 XN1 nS 0 intN1 RV523_NMOS
 XN2 nQ intN1 Q RV523_NMOS
 XN3 nR 0 intN2 RV523_NMOS
 XN4 Q intN2 nQ RV523_NMOS
 XP1 nS VDD Q RV523_PMOS
 XP2 nQ VDD Q RV523_PMOS
 XP3 nR VDD nQ RV523_PMOS
 XP4 Q VDD nQ RV523_PMOS
.ends
