VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

SITE CoreSite
  CLASS CORE ;
  SIZE 1 BY 4 ;
END CoreSite

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    SPACING 0.1 ;
    WIDTH 0.1 ;
    PITCH 0.2 ;
END M1
LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    SPACING 0.1 ;
    WIDTH 0.1 ;
    PITCH 0.2 ;
END M2

MACRO DECAP
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 1 BY 4 ;
  SITE CoreSite ;
END DECAP

MACRO DECAP_LED
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2 BY 4 ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 1.1 0.55 1.5 0.95 ;
    END
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 1.1 3.05 1.5 3.45 ;
    END
  END Y
END DECAP_LED

MACRO NOT
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 2 BY 4 ;
  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 1.3 1.55 1.7 1.95 ;
    END
  END Y
END NOT

MACRO NAND2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4 BY 4 ;
  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 3.3 1.55 3.7 1.95 ;
    END
  END Y
END NAND2


MACRO NAND3
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 6 BY 4 ;
  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 5.3 1.55 5.7 1.95 ;
    END
  END Y
END NAND3

MACRO NAND4
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 8 BY 4 ;
  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 6.3 2.05 6.7 2.45 ;
    END
  END A4

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 7.3 1.55 7.7 1.95 ;
    END
  END Y
END NAND4

MACRO NOR2
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 4 BY 4 ;
  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 3.3 1.55 3.7 1.95 ;
    END
  END Y
END NOR2

MACRO NOR3
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 6 BY 4 ;
  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END A3

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 5.3 1.55 5.7 1.95 ;
    END
  END Y
END NOR3

MACRO NOR4
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 8 BY 4 ;
  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 6.3 2.05 6.7 2.45 ;
    END
  END A4

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 7.3 1.55 7.7 1.95 ;
    END
  END Y
END NOR4

MACRO AOI22
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 8 BY 4 ;

  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 6.3 2.05 6.7 2.45 ;
    END
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 7.3 1.55 7.7 1.95 ;
    END
  END Y

END AOI22

MACRO OAI22
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 8 BY 4 ;

  SITE CoreSite ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 6.3 2.05 6.7 2.45 ;
    END
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 7.3 1.55 7.7 1.95 ;
    END
  END Y

END OAI22

MACRO AOI211
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 8 BY 4 ;

  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 6.3 2.05 6.7 2.45 ;
    END
  END C2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 7.3 1.55 7.7 1.95 ;
    END
  END Y

END AOI211

MACRO OAI211
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 8 BY 4 ;

  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 6.3 2.05 6.7 2.45 ;
    END
  END C2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 7.3 1.55 7.7 1.95 ;
    END
  END Y

END OAI211

MACRO AOI21
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 6 BY 4 ;

  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 5.3 1.55 5.7 2.45 ;
    END
  END Y

END AOI21


MACRO OAI21
  CLASS CORE ;
  ORIGIN 0 0 ;
  SIZE 6 BY 4 ;

  SITE CoreSite ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 0.3 2.05 0.7 2.45 ;
    END
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 2.3 2.05 2.7 2.45 ;
    END
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 4.3 2.05 4.7 2.45 ;
    END
  END B2

  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
      RECT 5.3 1.55 5.7 1.95 ;
    END
  END Y

END OAI21


END LIBRARY