* Main ngspice simulation file

.include "OAI22.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A1 A2 B1 B2 OAI22

.TRAN 0.1ns 48200ns

* Simulation control
.control 
    run
    write OAI22.raw
    quit
.endc
.END