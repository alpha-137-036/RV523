* Main ngspice simulation file

.include "AOI21.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A B1 B2 AOI21

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write AOI21.raw
    quit
.endc
.END