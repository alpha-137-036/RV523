* Main ngspice simulation file

.include "D_FLIP_FLOP.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on outputs
CloadQ Q 0 30p
CloadnQ nQ 0 30p

* Instantiate D_FLIP_FLOP gate
XU1 Q nQ D EN nEN D_FLIP_FLOP

.TRAN 0.1ns 1200ns

* Simulation control
.control 
    run
    write D_FLIP_FLOP.raw
    quit
.endc
.END