.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt NAND2 Y A1 A2
 XN1 A1 0 int1 RV523_NMOS
 XN2 A2 int1 Y RV523_NMOS
 XP1 A1 VDD Y RV523_PMOS
 XP2 A2 VDD Y RV523_PMOS
.ends
