* Main ngspice simulation file

.include "../RV523_global.sp"
.include "NOT.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate cell
XU1 Y A VDD 0 NOT

.TRAN 0.1ns 600ns

* Simulation control
.control 
    run
    write NOT.raw
    quit
.endc
.END