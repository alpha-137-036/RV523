* Main ngspice simulation file

.include "../RV523_global.sp"
.include "AOI211.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A B C1 C2 VDD 0 AOI211

.TRAN 0.1ns 48200ns

* Simulation control
.control 
    run
    write AOI211.raw
    quit
.endc
.END