.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt NOT Y A
 XN1 A 0 Y RV523_NMOS
 XP1 A VDD Y RV523_PMOS
.ends
