.subckt AOI22 Y A1 A2 B1 B2 VDD VSS
 XN1 A1 VSS intA RV523_NMOS
 XN2 A2 intA Y RV523_NMOS
 XN3 B1 VSS intB RV523_NMOS
 XN4 B2 intB Y RV523_NMOS
 XP1 A1 intP Y RV523_PMOS
 XP2 A2 intP Y RV523_PMOS
 XP3 B1 VDD intP RV523_PMOS
 XP4 B2 VDD intP RV523_PMOS
.ends
