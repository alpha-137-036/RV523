.model G2N7002X_CORE NMOS (VTO=1.40 KP=5.25e-08 L=5.26e-04 W=1.45e-02)
.model SP2006KT5_CORE PMOS (VTO=-0.65 KP=3.568e-06 W=1 L=3.053e-05)

* G2N7002X NMOS Subcircuit
.subckt G2N7002X D G S B
* Internal node for drain after Rds(on)
X1 D_INT G S B G2N7002X_CORE
RDS D D_INT 1.3
Cgs G S 33p
Cgd G D_INT 17p
.ends G2N7002X

* SP2006KT5 PMOS Subcircuit
.subckt SP2006KT5 D G S B
* Internal node for drain after Rds(on)
X1 D_INT G S B SP2006KT5_CORE
RDS D D_INT 0.85
Cgs G S 75p
Cgd G D_INT 38p
.ends SP2006KT5

* Inverter using G2N7002X and SP2006KT5
VDD VDD 0 DC 1.8
VIN IN 0 PULSE(0 1.8 0 1n 1n 500n 1u)
X1 OUT IN 0 0 G2N7002X
X2 OUT IN VDD VDD SP2006KT5
CL OUT 0 5p

* Simulation control
.tran 1n 2u
.control
run
plot VIN OUT
.endc

.end

