(* blackbox *)
(* footprint="Package_TO_SOT_SMD:SOT-523" *)
module NMOS(
    (* num="1" *)
    inout G, 
    (* num="3" *)
    inout D,
    (* num="2" *)
    inout S
);
endmodule

(* blackbox *)
(* footprint="Package_TO_SOT_SMD:SOT-523" *)
module PMOS(
    (* num="1" *)
    inout G, 
    (* num="3" *)
    inout D,
    (* num="2" *)
    inout S
);
endmodule

