* Main ngspice simulation file

.include "NAND.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate NAND gate
XU1 Y A B NAND

.TRAN 0.1ns 2600ns

* Simulation control
.control 
    run
    write NAND.raw
    quit
.endc
.END