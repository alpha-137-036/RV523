* Main ngspice simulation file

.include "NOR.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate NOR gate
XU1 Y A B NOR

.TRAN 0.1ns 2600ns

* Simulation control
.control 
    run
    write NOR.raw
    quit
.endc
.END