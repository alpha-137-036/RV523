* Main ngspice simulation file

.include "NOR2.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate NOR2 gate
XU1 Y A1 A2 NOR2

.TRAN 0.1ns 2600ns

* Simulation control
.control 
    run
    write NOR2.raw
    quit
.endc
.END