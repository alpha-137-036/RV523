* Main ngspice simulation file

.include "../RV523_global.sp"
.include "NOR4.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate cell
XU1 Y A1 A2 A3 A4 VDD 0 NOR4

.TRAN 0.1ns 49000ns

* Simulation control
.control 
    run
    write NOR4.raw
    quit
.endc
.END