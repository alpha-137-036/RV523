.subckt OR3 Y A1 A2 A3 VDD VSS
 Xnor1.N1 A1 VSS nY RV523_NMOS
 Xnor1.N2 A2 VSS nY RV523_NMOS
 Xnor1.N3 A3 VSS nY RV523_NMOS
 Xnor1.P1 A1 nor1.int1 nY RV523_PMOS
 Xnor1.P2 A2 nor1.int2 nor1.int1 RV523_PMOS
 Xnor1.P3 A3 VDD nor1.int2 RV523_PMOS
 Xnot1.N1 nY VSS Y RV523_NMOS
 Xnot1.P1 nY VDD Y RV523_PMOS
.ends
