.subckt D_LATCH Q nQ D CLK nCLK VDD VSS
 XNOT1.N1 D VSS NOT1.intN RV523_NMOS
 XNOT1.N2 CLK NOT1.intN nQ RV523_NMOS
 XNOT1.P1 D VDD NOT1.intP RV523_PMOS
 XNOT1.P2 nCLK NOT1.intP nQ RV523_PMOS
 XNOT2.N1 nQ VSS Q RV523_NMOS
 XNOT2.P1 nQ VDD Q RV523_PMOS
 XNOT3.N1 Q VSS NOT3.intN RV523_NMOS
 XNOT3.N2 nCLK NOT3.intN nQ RV523_NMOS
 XNOT3.P1 Q VDD NOT3.intP RV523_PMOS
 XNOT3.P2 CLK NOT3.intP nQ RV523_PMOS
.ends
