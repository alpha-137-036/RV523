module DECAP_LED(
    input A,
    input LED_GND
);
endmodule