.subckt NAND4 Y A1 A2 A3 A4 VDD VSS
 XN1 A1 VSS int1 RV523_NMOS
 XN2 A2 int1 int2 RV523_NMOS
 XN3 A3 int2 int3 RV523_NMOS
 XN4 A4 int3 Y RV523_NMOS
 XP1 A1 VDD Y RV523_PMOS
 XP2 A2 VDD Y RV523_PMOS
 XP3 A3 VDD Y RV523_PMOS
 XP4 A4 VDD Y RV523_PMOS
.ends
