.subckt TINV Y A EN nEN VDD VSS
 XN1 A VSS intN RV523_NMOS
 XN2 EN intN Y RV523_NMOS
 XP1 A VDD intP RV523_PMOS
 XP2 nEN intP Y RV523_PMOS
.ends
