* Main ngspice simulation file

.include "../RV523_global.sp"
.include "NAND2.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate NAND gate
XU1 Y A1 A2 VDD 0 NAND2

.TRAN 0.1ns 2600ns

* Simulation control
.control 
    run
    write NAND2.raw
    quit
.endc
.END