* Main ngspice simulation file

.include "NAND4.ckt"
.include "pwl_Inputs.sp"

.global VDD

.ic V(Y)=0


VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate NAND4 gate
XU1 Y A1 A2 A3 A4 NAND4

.options abstol=1n vabstol=1u iabstol=1p reltol=1e-4
.TRAN 0.1ns 49000ns

* Simulation control
.control 
    run
    write NAND4.raw
    quit
.endc
.END