VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

SITE CoreSite
  CLASS CORE ;
  SIZE 1 BY 4 ;
END CoreSite

LAYER M1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    SPACING 0.1 ;
    WIDTH 0.1 ;
    PITCH 0.2 ;
END M1
LAYER M2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    SPACING 0.1 ;
    WIDTH 0.1 ;
    PITCH 0.2 ;
END M2


END LIBRARY