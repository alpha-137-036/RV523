.subckt OAI21 Y A B1 B2 VDD VSS
 XN1 A VSS intN RV523_NMOS
 XN2 B1 intN Y RV523_NMOS
 XN3 B2 intN Y RV523_NMOS
 XP1 A VDD Y RV523_PMOS
 XP2 B1 VDD intB RV523_PMOS
 XP3 B2 intB Y RV523_PMOS
.ends
