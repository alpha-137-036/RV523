* Main ngspice simulation file

.include "../RV523_global.sp"
.include "D_LATCH.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on outputs
CloadQ Q 0 30p
CloadnQ nQ 0 30p

* Instantiate D_LATCH gate
XU1 Q nQ D CLK nCLK VDD 0 D_LATCH

.TRAN 0.1ns 1200ns

* Simulation control
.control 
    run
    write D_LATCH.raw
    quit
.endc
.END