* Main ngspice simulation file

.include "NOT.ckt"
.include "pwl_Inputs.sp"
.include "../2n7002.sub"
.include "../bss84.sub"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate cell
XU1 A Y NOT

.TRAN 0.1ns 600ns

* Simulation control
.control 
    run
    write NOT.raw
    quit
.endc
.END