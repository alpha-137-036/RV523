* Main ngspice simulation file

.include "AOI211.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A B C1 C2 AOI211

.TRAN 0.1ns 48200ns

* Simulation control
.control 
    run
    write AOI211.raw
    quit
.endc
.END