* Main ngspice simulation file

.include "../RV523_global.sp"
.include "AOI22.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A1 A2 B1 B2 VDD 0 AOI22

.TRAN 0.1ns 48200ns

* Simulation control
.control 
    run
    write AOI22.raw
    quit
.endc
.END