* Main ngspice simulation file

.include "NOT.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate cell
XU1 Y A NOT

.TRAN 0.1ns 600ns

* Simulation control
.control 
    run
    write NOT.raw
    quit
.endc
.END