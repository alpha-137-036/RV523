.inc "2n7002.sub"
* SOT-523 pin order 1=G, 2=D, 3=S
.SUBCKT RV523_NMOS G S D
    * 2n7002 model has pin order D  G  S
    X1 D G S N7002
.ENDS
