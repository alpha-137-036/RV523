* Main ngspice simulation file

.include "NAND3.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 3.3

* Load capacitor on output
Cload Y 0 30p

* Instantiate NAND gate
XU1 Y A1 A2 A3 NAND3

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write NAND3.raw
    quit
.endc
.END