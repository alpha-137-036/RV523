.inc "RV523_NMOS.ckt"
.inc "RV523_PMOS.ckt"

.PARAM vdd=5V