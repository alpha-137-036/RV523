* Main ngspice simulation file

.inc "../RV523_global.sp"
.include "AOI21.ckt"
.include "pwl_Inputs.sp"

VDD VDD 0 {vdd}

* Load capacitor on output
Cload Y 0 30p

* Instantiate gate
XU1 Y A B1 B2 VDD 0 AOI21

.TRAN 0.1ns 11400ns

* Simulation control
.control 
    run
    write AOI21.raw
    quit
.endc
.END