* Main ngspice simulation file

.include "NOR4.ckt"
.include "pwl_Inputs.sp"

.global VDD

VDD VDD 0 5

* Load capacitor on output
Cload Y 0 30p

* Instantiate cell
XU1 Y A1 A2 A3 A4 NOR4

.TRAN 0.1ns 49000ns

* Simulation control
.control 
    run
    write NOR4.raw
    quit
.endc
.END