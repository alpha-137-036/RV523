(* blackbox *)
(* footprint="RV523:SOT523" *)
(* value="NMOS" *)
module RV523_NMOS(
    (* num="3" *)
    inout D,
    (* num="1" *)
    inout G, 
    (* num="2" *)
    inout S
);
endmodule

(* blackbox *)
(* footprint="RV523:SOT523" *)
(* value="PMOS" *)
module RV523_PMOS(
    (* num="3" *)
    inout D,
    (* num="1" *)
    inout G, 
    (* num="2" *)
    inout S
);
endmodule

