.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt AOI21 Y A B1 B2
 XN1 A 0 Y RV523_NMOS
 XN2 B1 0 intB RV523_NMOS
 XN3 B2 intB Y RV523_NMOS
 XP1 A intP Y RV523_PMOS
 XP2 B1 VDD intP RV523_PMOS
 XP3 B2 VDD intP RV523_PMOS
.ends
