.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt OAI211 Y A B C1 C2
 XN1 A 0 intNA RV523_NMOS
 XN2 B intNA intNB RV523_NMOS
 XN3 C1 intNB Y RV523_NMOS
 XN4 C2 intNB Y RV523_NMOS
 XP1 A VDD Y RV523_PMOS
 XP2 B VDD Y RV523_PMOS
 XP3 C1 VDD intC RV523_PMOS
 XP4 C2 intC Y RV523_PMOS
.ends
