.inc "../RV523_NMOS.ckt"
.inc "../RV523_PMOS.ckt"
.subckt NAND3 Y A B C
 XN1 A 0 int1 RV523_NMOS
 XN2 B int1 int2 RV523_NMOS
 XN3 C int2 Y RV523_NMOS
 XP1 A VDD Y RV523_PMOS
 XP2 B VDD Y RV523_PMOS
 XP3 C VDD Y RV523_PMOS
.ends
